** sch_path: /mnt/c/Users/NITHIN P/tb_opamp1.sch
**.subckt tb_opamp1
x2 START_N START VCC VSS not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=1
V2 VCC VSS 1.8
x4 ADJ DIFFOUT_N START START_N VCC VSS passgate W_N=0.5 L_N=0.15 W_P=0.5 L_P=0.15 m=1
XC2 ADJ VSS sky130_fd_pr__cap_mim_m3_2 W=10 L=10 MF=5 m=5
x5 DIFFOUT_N PLUS MINUS EN_N ADJ VCC VSS opam
**** begin user architecture code

.param mc_mm_switch=1
.param mc_pr_switch=0
.include /home/nithinpuru/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/nithinpuru/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/nithinpuru/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/nithinpuru/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice


* .option SCALE=1e-6
.option method=gear

* this experimental option enables mos model bin
* selection based on W/NF instead of W
.option wnflag=1


.param VCCGAUSS = agauss(1.8, 0.05, 1)
.param VCC = VCCGAUSS
** use of following line to remove VCC variations
* .param VCC =1.8

.param TEMPGAUSS = agauss(40, 30, 1)
.option temp = TEMPGAUSS
** use of following line to remove temperature variations
* .option temp =25

.include stimuli_tb_opamp.cir
.control
 option seed=9
 let run=0
 dowhile run <= 100
   save all
   tran 1n 4000n uic
   remzerovec
   write tb_opamp.raw
   set appendwrite
   reset
   let run = run + 1
 end
.endc




















**** end user architecture code
**.ends

* expanding   symbol:  sky130_tests/not.sym # of pins=2
** sym_path: /home/nithinpuru/pdk/sky130A/libs.tech/xschem/sky130_tests/not.sym
** sch_path: /home/nithinpuru/pdk/sky130A/libs.tech/xschem/sky130_tests/not.sch
.subckt not y a VCCPIN VSSPIN     W_N=1 L_N=0.15 W_P=2 L_P=0.15
*.opin y
*.ipin a
XM1 y a VSSPIN VSSPIN sky130_fd_pr__nfet_01v8 L=L_N W=W_N nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 y a VCCPIN VCCPIN sky130_fd_pr__pfet_01v8 L=L_P W=W_P nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  sky130_tests/passgate.sym # of pins=4
** sym_path: /home/nithinpuru/pdk/sky130A/libs.tech/xschem/sky130_tests/passgate.sym
** sch_path: /home/nithinpuru/pdk/sky130A/libs.tech/xschem/sky130_tests/passgate.sch
.subckt passgate Z A GP GN VCCBPIN VSSBPIN  W_N=1 L_N=0.2 W_P=1 L_P=0.2
*.iopin A
*.iopin Z
*.ipin GP
*.ipin GN
XM1 Z GN A VSSBPIN sky130_fd_pr__nfet_01v8 L=L_N W=W_N nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Z GP A VCCBPIN sky130_fd_pr__pfet_01v8 L=L_P W=W_P nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
* noconn VCCBPIN
* noconn VSSBPIN
.ends


* expanding   symbol:  /mnt/c/Users/NITHIN P/opam.sym # of pins=7
** sym_path: /mnt/c/Users/NITHIN P/opam.sym
** sch_path: /mnt/c/Users/NITHIN P/opam.sch
.subckt opam DIFFOUT_N PLUS MINUS EN_N ADJ VCC VSS
.ends

.end
