** sch_path: /home/nithinpuru/pdk/sky130A/libs.tech/xschem/sky130_tests/zero_opamp.sch
.subckt zero_opamp EN_N MINUS PLUS DIFFOUT VCC VSS ADJ
*.PININFO PLUS:I MINUS:I EN_N:I VSS:I VCC:I DIFFOUT:O ADJ:I
C6 G1 0 2f m=1
XM4 net9 EN_N VCC VCC sky130_fd_pr__pfet_01v8 L=8 W=2 nf=1 m=1
XM18 G2 G2 net7 VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 m=1
XM2 G1 G1 net8 VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 m=1
XM20 G2 PLUS net10 VCC sky130_fd_pr__pfet_01v8_lvt L=2 W=8 nf=1 m=1
XM3 G1 MINUS net11 VCC sky130_fd_pr__pfet_01v8_lvt L=2 W=8 nf=1 m=1
v1 SP net11 0
.save i(v1)
C4 SP 0 2f m=1
C1 G2 0 2f m=1
C5 DIFFOUT 0 4f m=1
XM6 DIFFOUT G2 net1 VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 m=1
v2 SP net10 0
.save i(v2)
v4 net1 VSS 0
.save i(v4)
v6 net9 SP 0
.save i(v6)
XM7 DIFFOUT EN_N VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=1
XM46 net12 EN_N VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=5 nf=1 m=1
v17 net12 net3 0
.save i(v17)
XM12 net2 G1 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 m=1
XM54 net2 net2 net3 VCC sky130_fd_pr__pfet_01v8_lvt L=4 W=4 nf=1 m=1
XM5 DIFFOUT net2 net3 VCC sky130_fd_pr__pfet_01v8_lvt L=4 W=4 nf=1 m=1
XM8 net5 ADJ net4 VCC sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XM9 net5 ADJ net6 VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=0.5 nf=1 m=1
XM10 net6 VCC VSS VSS sky130_fd_pr__nfet_01v8_lvt L=8 W=0.5 nf=1 m=1
XM1 net4 EN_N VCC VCC sky130_fd_pr__pfet_01v8 L=8 W=1 nf=1 m=1
v3 net5 G1 0
.save i(v3)
v5 net7 VSS 0
.save i(v5)
v7 net8 VSS 0
.save i(v7)
.ends
.end
